always @ (posedge i_Clk)
begin
    and_gate <= input_1 & input_2;
end