process (input_1, input_2)
begin
    and_gate <= input_1 and input_2;
end